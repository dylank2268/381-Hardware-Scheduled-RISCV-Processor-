--Micahel Berg and Dylan Kramer 
--all 4 pipeline register test bench 